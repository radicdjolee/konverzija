----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/18/2023 07:33:48 AM
-- Design Name: 
-- Module Name: cos_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cos_rom is
    generic (
	       WIDTH : integer := 32;
	       WIDTH_2 : integer := 64;
	       WIDTH_3 : integer := 96; 
	       WADDR   : integer := 10
    );
    port(
        address_cos_0 : in  std_logic_vector(WADDR-1 downto 0);
        dout_cos_0    : out std_logic_vector(WIDTH-1 downto 0)
    );
end cos_rom;

architecture Behavioral of cos_rom is
  type mem is array ( 0 to 647) of std_logic_vector(WIDTH-1 downto 0);
  constant my_Rom : mem := (

0 => "00001010110011110011011101110110",
1 => "11110011010011100110110100010110",
2 => "11110111011001110011100000011101",
3 => "00001110001100010011001001110010",
4 => "00000110000111110111100000110110",
5 => "11110000101111011001001100111110",
6 => "11111100100010010111011000110110",
7 => "00001111110111001111010101101111",
8 => "00000000101100101010101001000010",
9 => "11110000000000111110011000111111",
10 => "00000010000101101010001001101110",
11 => "00001111100111101110100010001110",
12 => "11111011001100000100111011101000",
13 => "11110001001101111100100110011011",
14 => "00000111011000110101001011101011",
15 => "00001101011111101000011110010000",
16 => "11110110010000101000001111010011",
17 => "11110100001101000001110100001000",
18 => "00001001101111010111110000101101",
19 => "11110001001101111100100110011011",
20 => "11111101111010010101110110010010",
21 => "00001111110111001111010101101111",
22 => "11111001111000001000011111001010",
23 => "11110011010011100110110100010110",
24 => "00001100101100011001001011101010",
25 => "00000110000111110111100000110110",
26 => "11110000001000110000101010010001",
27 => "00000010000101101010001001101110",
28 => "00001110110010000011011001100101",
29 => "11110110010000101000001111010011",
30 => "11110110010000101000001111010011",
31 => "00001110110010000011011001100101",
32 => "00000010000101101010001001101110",
33 => "11110000001000110000101010010001",
34 => "00000110000111110111100000110110",
35 => "00001100101100011001001011101010",
36 => "00001000100110001100011111100011",
37 => "11110000001000110000101010010001",
38 => "00000100110011111011000100011000",
39 => "00001011110010111110001011111000",
40 => "11110001001101111100100110011011",
41 => "00000000101100101010101001000010",
42 => "00001110001100010011001001110010",
43 => "11110011010011100110110100010110",
44 => "11111100100010010111011000110110",
45 => "00001111100111101110100010001110",
46 => "11110110010000101000001111010011",
47 => "11111000100111001010110100010101",
48 => "00001111111111000001100111000001",
49 => "11111001111000001000011111001010",
50 => "11110101001100001100100010001010",
51 => "00001111010000100110110011000010",
52 => "11111101111010010101110110010010",
53 => "11110010100000010111100001110000",
54 => "00000111011000110101001011101011",
55 => "11110000001000110000101010010001",
56 => "00001010110011110011011101110110",
57 => "00000011011101101000100111001010",
58 => "11110001001101111100100110011011",
59 => "00001101011111101000011110010000",
60 => "11111111010011010101010110111110",
61 => "11110011010011100110110100010110",
62 => "00001111010000100110110011000010",
63 => "11111011001100000100111011101000",
64 => "11110110010000101000001111010011",
65 => "00001111111111000001100111000001",
66 => "11110111011001110011100000011101",
67 => "11111001111000001000011111001010",
68 => "00001111100111101110100010001110",
69 => "11110100001101000001110100001000",
70 => "11111101111010010101110110010010",
71 => "00001110001100010011001001110010",
72 => "00000110000111110111100000110110",
73 => "11110001001101111100100110011011",
74 => "00001110110010000011011001100101",
75 => "11111001111000001000011111001010",
76 => "11111001111000001000011111001010",
77 => "00001110110010000011011001100101",
78 => "11110001001101111100100110011011",
79 => "00000110000111110111100000110110",
80 => "00000110000111110111100000110110",
81 => "11110001001101111100100110011011",
82 => "00001110110010000011011001100101",
83 => "11111001111000001000011111001010",
84 => "11111001111000001000011111001010",
85 => "00001110110010000011011001100101",
86 => "11110001001101111100100110011011",
87 => "00000110000111110111100000110110",
88 => "00000110000111110111100000110110",
89 => "11110001001101111100100110011011",
90 => "00000100110011111011000100011000",
91 => "11110011010011100110110100010110",
92 => "00001111111111000001100111000001",
93 => "11110010100000010111100001110000",
94 => "00000110000111110111100000110110",
95 => "00000011011101101000100111001010",
96 => "11110100001101000001110100001000",
97 => "00001111110111001111010101101111",
98 => "11110001110011101100110110001110",
99 => "00000111011000110101001011101011",
100 => "00000010000101101010001001101110",
101 => "11110101001100001100100010001010",
102 => "00001111100111101110100010001110",
103 => "11110001001101111100100110011011",
104 => "00001000100110001100011111100011",
105 => "00000000101100101010101001000010",
106 => "11110110010000101000001111010011",
107 => "00001111010000100110110011000010",
108 => "00000011011101101000100111001010",
109 => "11110110010000101000001111010011",
110 => "00001110001100010011001001110010",
111 => "11110000000000111110011000111111",
112 => "00001110110010000011011001100101",
113 => "11110101001100001100100010001010",
114 => "00000100110011111011000100011000",
115 => "00000010000101101010001001101110",
116 => "11110111011001110011100000011101",
117 => "00001101011111101000011110010000",
118 => "11110000001000110000101010010001",
119 => "00001111010000100110110011000010",
120 => "11110100001101000001110100001000",
121 => "00000110000111110111100000110110",
122 => "00000000101100101010101001000010",
123 => "11111000100111001010110100010101",
124 => "00001100101100011001001011101010",
125 => "11110000011000010001011101110010",
126 => "00000010000101101010001001101110",
127 => "11111001111000001000011111001010",
128 => "00001001101111010111110000101101",
129 => "11110011010011100110110100010110",
130 => "00001110110010000011011001100101",
131 => "11110000001000110000101010010001",
132 => "00001111110111001111010101101111",
133 => "11110001001101111100100110011011",
134 => "00001100101100011001001011101010",
135 => "11110110010000101000001111010011",
136 => "00000110000111110111100000110110",
137 => "11111101111010010101110110010010",
138 => "11111101111010010101110110010010",
139 => "00000110000111110111100000110110",
140 => "11110110010000101000001111010011",
141 => "00001100101100011001001011101010",
142 => "11110001001101111100100110011011",
143 => "00001111110111001111010101101111",
144 => "00000000101100101010101001000010",
145 => "11111101111010010101110110010010",
146 => "00000011011101101000100111001010",
147 => "11111011001100000100111011101000",
148 => "00000110000111110111100000110110",
149 => "11111000100111001010110100010101",
150 => "00001000100110001100011111100011",
151 => "11110110010000101000001111010011",
152 => "00001010110011110011011101110110",
153 => "11110100001101000001110100001000",
154 => "00001100101100011001001011101010",
155 => "11110010100000010111100001110000",
156 => "00001110001100010011001001110010",
157 => "11110001001101111100100110011011",
158 => "00001111010000100110110011000010",
159 => "11110000011000010001011101110010",
160 => "00001111110111001111010101101111",
161 => "11110000000000111110011000111111",
162 => "11111111010011010101010110111110",
163 => "00000010000101101010001001101110",
164 => "11111100100010010111011000110110",
165 => "00000100110011111011000100011000",
166 => "11111001111000001000011111001010",
167 => "00000111011000110101001011101011",
168 => "11110111011001110011100000011101",
169 => "00001001101111010111110000101101",
170 => "11110101001100001100100010001010",
171 => "00001011110010111110001011111000",
172 => "11110011010011100110110100010110",
173 => "00001101011111101000011110010000",
174 => "11110001110011101100110110001110",
175 => "00001110110010000011011001100101",
176 => "11110000101111011001001100111110",
177 => "00001111100111101110100010001110",
178 => "11110000001000110000101010010001",
179 => "00001111111111000001100111000001",
180 => "11111101111010010101110110010010",
181 => "00000110000111110111100000110110",
182 => "11110110010000101000001111010011",
183 => "00001100101100011001001011101010",
184 => "11110001001101111100100110011011",
185 => "00001111110111001111010101101111",
186 => "11110000001000110000101010010001",
187 => "00001110110010000011011001100101",
188 => "11110011010011100110110100010110",
189 => "00001001101111010111110000101101",
190 => "11111001111000001000011111001010",
191 => "00000010000101101010001001101110",
192 => "00000010000101101010001001101110",
193 => "11111001111000001000011111001010",
194 => "00001001101111010111110000101101",
195 => "11110011010011100110110100010110",
196 => "00001110110010000011011001100101",
197 => "11110000001000110000101010010001",
198 => "11111100100010010111011000110110",
199 => "00001001101111010111110000101101",
200 => "11110001110011101100110110001110",
201 => "00001111111111000001100111000001",
202 => "11110001001101111100100110011011",
203 => "00001010110011110011011101110110",
204 => "11111011001100000100111011101000",
205 => "11111101111010010101110110010010",
206 => "00001000100110001100011111100011",
207 => "11110010100000010111100001110000",
208 => "00001111110111001111010101101111",
209 => "11110000101111011001001100111110",
210 => "00001011110010111110001011111000",
211 => "11111001111000001000011111001010",
212 => "11111111010011010101010110111110",
213 => "00000111011000110101001011101011",
214 => "11110011010011100110110100010110",
215 => "00001111100111101110100010001110",
216 => "11111011001100000100111011101000",
217 => "00001100101100011001001011101010",
218 => "11110000000000111110011000111111",
219 => "00001101011111101000011110010000",
220 => "11111001111000001000011111001010",
221 => "11111100100010010111011000110110",
222 => "00001011110010111110001011111000",
223 => "11110000001000110000101010010001",
224 => "00001110001100010011001001110010",
225 => "11111000100111001010110100010101",
226 => "11111101111010010101110110010010",
227 => "00001010110011110011011101110110",
228 => "11110000011000010001011101110010",
229 => "00001110110010000011011001100101",
230 => "11110111011001110011100000011101",
231 => "11111111010011010101010110111110",
232 => "00001001101111010111110000101101",
233 => "11110000101111011001001100111110",
234 => "11111001111000001000011111001010",
235 => "00001110110010000011011001100101",
236 => "11110001001101111100100110011011",
237 => "00000110000111110111100000110110",
238 => "00000110000111110111100000110110",
239 => "11110001001101111100100110011011",
240 => "00001110110010000011011001100101",
241 => "11111001111000001000011111001010",
242 => "11111001111000001000011111001010",
243 => "00001110110010000011011001100101",
244 => "11110001001101111100100110011011",
245 => "00000110000111110111100000110110",
246 => "00000110000111110111100000110110",
247 => "11110001001101111100100110011011",
248 => "00001110110010000011011001100101",
249 => "11111001111000001000011111001010",
250 => "11111001111000001000011111001010",
251 => "00001110110010000011011001100101",
252 => "11111000100111001010110100010101",
253 => "00001111110111001111010101101111",
254 => "11110101001100001100100010001010",
255 => "11111100100010010111011000110110",
256 => "00001110110010000011011001100101",
257 => "11110010100000010111100001110000",
258 => "00000000101100101010101001000010",
259 => "00001100101100011001001011101010",
260 => "11110000101111011001001100111110",
261 => "00000100110011111011000100011000",
262 => "00001001101111010111110000101101",
263 => "11110000000000111110011000111111",
264 => "00001000100110001100011111100011",
265 => "00000110000111110111100000110110",
266 => "11110000011000010001011101110010",
267 => "00001011110010111110001011111000",
268 => "00000010000101101010001001101110",
269 => "11110001110011101100110110001110",
270 => "11110111011001110011100000011101",
271 => "00001111110111001111010101101111",
272 => "11111011001100000100111011101000",
273 => "11110100001101000001110100001000",
274 => "00001110110010000011011001100101",
275 => "11111111010011010101010110111110",
276 => "11110001110011101100110110001110",
277 => "00001100101100011001001011101010",
278 => "00000011011101101000100111001010",
279 => "11110000011000010001011101110010",
280 => "00001001101111010111110000101101",
281 => "00000111011000110101001011101011",
282 => "11110000000000111110011000111111",
283 => "00000110000111110111100000110110",
284 => "00001010110011110011011101110110",
285 => "11110000101111011001001100111110",
286 => "00000010000101101010001001101110",
287 => "00001101011111101000011110010000",
288 => "11110110010000101000001111010011",
289 => "00001110110010000011011001100101",
290 => "00000010000101101010001001101110",
291 => "11110000001000110000101010010001",
292 => "00000110000111110111100000110110",
293 => "00001100101100011001001011101010",
294 => "11110011010011100110110100010110",
295 => "11111001111000001000011111001010",
296 => "00001111110111001111010101101111",
297 => "11111101111010010101110110010010",
298 => "11110001001101111100100110011011",
299 => "00001001101111010111110000101101",
300 => "00001001101111010111110000101101",
301 => "11110001001101111100100110011011",
302 => "11111101111010010101110110010010",
303 => "00001111110111001111010101101111",
304 => "11111001111000001000011111001010",
305 => "11110011010011100110110100010110",
306 => "11110101001100001100100010001010",
307 => "00001100101100011001001011101010",
308 => "00001000100110001100011111100011",
309 => "11110001110011101100110110001110",
310 => "11111001111000001000011111001010",
311 => "00001111010000100110110011000010",
312 => "00000011011101101000100111001010",
313 => "11110000001000110000101010010001",
314 => "11111111010011010101010110111110",
315 => "00001111111111000001100111000001",
316 => "11111101111010010101110110010010",
317 => "11110000011000010001011101110010",
318 => "00000100110011111011000100011000",
319 => "00001110110010000011011001100101",
320 => "11111000100111001010110100010101",
321 => "11110010100000010111100001110000",
322 => "00001001101111010111110000101101",
323 => "00001011110010111110001011111000",
324 => "11110100001101000001110100001000",
325 => "00001001101111010111110000101101",
326 => "00001101011111101000011110010000",
327 => "11111000100111001010110100010101",
328 => "11110001001101111100100110011011",
329 => "00000100110011111011000100011000",
330 => "00001111100111101110100010001110",
331 => "11111101111010010101110110010010",
332 => "11110000000000111110011000111111",
333 => "11111111010011010101010110111110",
334 => "00001111110111001111010101101111",
335 => "00000011011101101000100111001010",
336 => "11110000101111011001001100111110",
337 => "11111001111000001000011111001010",
338 => "00001110001100010011001001110010",
339 => "00001000100110001100011111100011",
340 => "11110011010011100110110100010110",
341 => "11110101001100001100100010001010",
342 => "11110011010011100110110100010110",
343 => "00000110000111110111100000110110",
344 => "00001111110111001111010101101111",
345 => "00000010000101101010001001101110",
346 => "11110001001101111100100110011011",
347 => "11110110010000101000001111010011",
348 => "00001001101111010111110000101101",
349 => "00001110110010000011011001100101",
350 => "11111101111010010101110110010010",
351 => "11110000001000110000101010010001",
352 => "11111001111000001000011111001010",
353 => "00001100101100011001001011101010",
354 => "00001100101100011001001011101010",
355 => "11111001111000001000011111001010",
356 => "11110000001000110000101010010001",
357 => "11111101111010010101110110010010",
358 => "00001110110010000011011001100101",
359 => "00001001101111010111110000101101",
360 => "11110010100000010111100001110000",
361 => "00000010000101101010001001101110",
362 => "00001111010000100110110011000010",
363 => "00001010110011110011011101110110",
364 => "11111001111000001000011111001010",
365 => "11110000000000111110011000111111",
366 => "11111000100111001010110100010101",
367 => "00001001101111010111110000101101",
368 => "00001111100111101110100010001110",
369 => "00000011011101101000100111001010",
370 => "11110011010011100110110100010110",
371 => "11110001110011101100110110001110",
372 => "00000000101100101010101001000010",
373 => "00001110110010000011011001100101",
374 => "00001011110010111110001011111000",
375 => "11111011001100000100111011101000",
376 => "11110000001000110000101010010001",
377 => "11110111011001110011100000011101",
378 => "11110001110011101100110110001110",
379 => "11111101111010010101110110010010",
380 => "00001011110010111110001011111000",
381 => "00001111100111101110100010001110",
382 => "00000110000111110111100000110110",
383 => "11110111011001110011100000011101",
384 => "11110000000000111110011000111111",
385 => "11110110010000101000001111010011",
386 => "00000100110011111011000100011000",
387 => "00001111010000100110110011000010",
388 => "00001100101100011001001011101010",
389 => "11111111010011010101010110111110",
390 => "11110010100000010111100001110000",
391 => "11110001001101111100100110011011",
392 => "11111100100010010111011000110110",
393 => "00001010110011110011011101110110",
394 => "00001111110111001111010101101111",
395 => "00000111011000110101001011101011",
396 => "11110001001101111100100110011011",
397 => "11111001111000001000011111001010",
398 => "00000110000111110111100000110110",
399 => "00001110110010000011011001100101",
400 => "00001110110010000011011001100101",
401 => "00000110000111110111100000110110",
402 => "11111001111000001000011111001010",
403 => "11110001001101111100100110011011",
404 => "11110001001101111100100110011011",
405 => "11111001111000001000011111001010",
406 => "00000110000111110111100000110110",
407 => "00001110110010000011011001100101",
408 => "00001110110010000011011001100101",
409 => "00000110000111110111100000110110",
410 => "11111001111000001000011111001010",
411 => "11110001001101111100100110011011",
412 => "11110001001101111100100110011011",
413 => "11111001111000001000011111001010",
414 => "11110000101111011001001100111110",
415 => "11110110010000101000001111010011",
416 => "11111111010011010101010110111110",
417 => "00001000100110001100011111100011",
418 => "00001110110010000011011001100101",
419 => "00001111100111101110100010001110",
420 => "00001010110011110011011101110110",
421 => "00000010000101101010001001101110",
422 => "11111000100111001010110100010101",
423 => "11110001110011101100110110001110",
424 => "11110000001000110000101010010001",
425 => "11110100001101000001110100001000",
426 => "11111100100010010111011000110110",
427 => "00000110000111110111100000110110",
428 => "00001101011111101000011110010000",
429 => "00001111111111000001100111000001",
430 => "00001100101100011001001011101010",
431 => "00000100110011111011000100011000",
432 => "11110000011000010001011101110010",
433 => "11110011010011100110110100010110",
434 => "11111000100111001010110100010101",
435 => "11111111010011010101010110111110",
436 => "00000110000111110111100000110110",
437 => "00001011110010111110001011111000",
438 => "00001111010000100110110011000010",
439 => "00001111110111001111010101101111",
440 => "00001101011111101000011110010000",
441 => "00001000100110001100011111100011",
442 => "00000010000101101010001001101110",
443 => "11111011001100000100111011101000",
444 => "11110101001100001100100010001010",
445 => "11110001001101111100100110011011",
446 => "11110000000000111110011000111111",
447 => "11110001110011101100110110001110",
448 => "11110110010000101000001111010011",
449 => "11111100100010010111011000110110",
450 => "11110000001000110000101010010001",
451 => "11110001001101111100100110011011",
452 => "11110011010011100110110100010110",
453 => "11110110010000101000001111010011",
454 => "11111001111000001000011111001010",
455 => "11111101111010010101110110010010",
456 => "00000010000101101010001001101110",
457 => "00000110000111110111100000110110",
458 => "00001001101111010111110000101101",
459 => "00001100101100011001001011101010",
460 => "00001110110010000011011001100101",
461 => "00001111110111001111010101101111",
462 => "00001111110111001111010101101111",
463 => "00001110110010000011011001100101",
464 => "00001100101100011001001011101010",
465 => "00001001101111010111110000101101",
466 => "00000110000111110111100000110110",
467 => "00000010000101101010001001101110",
468 => "11110000000000111110011000111111",
469 => "11110000001000110000101010010001",
470 => "11110000011000010001011101110010",
471 => "11110000101111011001001100111110",
472 => "11110001001101111100100110011011",
473 => "11110001110011101100110110001110",
474 => "11110010100000010111100001110000",
475 => "11110011010011100110110100010110",
476 => "11110100001101000001110100001000",
477 => "11110101001100001100100010001010",
478 => "11110110010000101000001111010011",
479 => "11110111011001110011100000011101",
480 => "11111000100111001010110100010101",
481 => "11111001111000001000011111001010",
482 => "11111011001100000100111011101000",
483 => "11111100100010010111011000110110",
484 => "11111101111010010101110110010010",
485 => "11111111010011010101010110111110",
486 => "11110000000000111110011000111111",
487 => "11110000001000110000101010010001",
488 => "11110000011000010001011101110010",
489 => "11110000101111011001001100111110",
490 => "11110001001101111100100110011011",
491 => "11110001110011101100110110001110",
492 => "11110010100000010111100001110000",
493 => "11110011010011100110110100010110",
494 => "11110100001101000001110100001000",
495 => "11110101001100001100100010001010",
496 => "11110110010000101000001111010011",
497 => "11110111011001110011100000011101",
498 => "11111000100111001010110100010101",
499 => "11111001111000001000011111001010",
500 => "11111011001100000100111011101000",
501 => "11111100100010010111011000110110",
502 => "11111101111010010101110110010010",
503 => "11111111010011010101010110111110",
504 => "11110000001000110000101010010001",
505 => "11110001001101111100100110011011",
506 => "11110011010011100110110100010110",
507 => "11110110010000101000001111010011",
508 => "11111001111000001000011111001010",
509 => "11111101111010010101110110010010",
510 => "00000010000101101010001001101110",
511 => "00000110000111110111100000110110",
512 => "00001001101111010111110000101101",
513 => "00001100101100011001001011101010",
514 => "00001110110010000011011001100101",
515 => "00001111110111001111010101101111",
516 => "00001111110111001111010101101111",
517 => "00001110110010000011011001100101",
518 => "00001100101100011001001011101010",
519 => "00001001101111010111110000101101",
520 => "00000110000111110111100000110110",
521 => "00000010000101101010001001101110",
522 => "11110000011000010001011101110010",
523 => "11110011010011100110110100010110",
524 => "11111000100111001010110100010101",
525 => "11111111010011010101010110111110",
526 => "00000110000111110111100000110110",
527 => "00001011110010111110001011111000",
528 => "00001111010000100110110011000010",
529 => "00001111110111001111010101101111",
530 => "00001101011111101000011110010000",
531 => "00001000100110001100011111100011",
532 => "00000010000101101010001001101110",
533 => "11111011001100000100111011101000",
534 => "11110101001100001100100010001010",
535 => "11110001001101111100100110011011",
536 => "11110000000000111110011000111111",
537 => "11110001110011101100110110001110",
538 => "11110110010000101000001111010011",
539 => "11111100100010010111011000110110",
540 => "11110000101111011001001100111110",
541 => "11110110010000101000001111010011",
542 => "11111111010011010101010110111110",
543 => "00001000100110001100011111100011",
544 => "00001110110010000011011001100101",
545 => "00001111100111101110100010001110",
546 => "00001010110011110011011101110110",
547 => "00000010000101101010001001101110",
548 => "11111000100111001010110100010101",
549 => "11110001110011101100110110001110",
550 => "11110000001000110000101010010001",
551 => "11110100001101000001110100001000",
552 => "11111100100010010111011000110110",
553 => "00000110000111110111100000110110",
554 => "00001101011111101000011110010000",
555 => "00001111111111000001100111000001",
556 => "00001100101100011001001011101010",
557 => "00000100110011111011000100011000",
558 => "11110001001101111100100110011011",
559 => "11111001111000001000011111001010",
560 => "00000110000111110111100000110110",
561 => "00001110110010000011011001100101",
562 => "00001110110010000011011001100101",
563 => "00000110000111110111100000110110",
564 => "11111001111000001000011111001010",
565 => "11110001001101111100100110011011",
566 => "11110001001101111100100110011011",
567 => "11111001111000001000011111001010",
568 => "00000110000111110111100000110110",
569 => "00001110110010000011011001100101",
570 => "00001110110010000011011001100101",
571 => "00000110000111110111100000110110",
572 => "11111001111000001000011111001010",
573 => "11110001001101111100100110011011",
574 => "11110001001101111100100110011011",
575 => "11111001111000001000011111001010",
576 => "11110001110011101100110110001110",
577 => "11111101111010010101110110010010",
578 => "00001011110010111110001011111000",
579 => "00001111100111101110100010001110",
580 => "00000110000111110111100000110110",
581 => "11110111011001110011100000011101",
582 => "11110000000000111110011000111111",
583 => "11110110010000101000001111010011",
584 => "00000100110011111011000100011000",
585 => "00001111010000100110110011000010",
586 => "00001100101100011001001011101010",
587 => "11111111010011010101010110111110",
588 => "11110010100000010111100001110000",
589 => "11110001001101111100100110011011",
590 => "11111100100010010111011000110110",
591 => "00001010110011110011011101110110",
592 => "00001111110111001111010101101111",
593 => "00000111011000110101001011101011",
594 => "11110010100000010111100001110000",
595 => "00000010000101101010001001101110",
596 => "00001111010000100110110011000010",
597 => "00001010110011110011011101110110",
598 => "11111001111000001000011111001010",
599 => "11110000000000111110011000111111",
600 => "11111000100111001010110100010101",
601 => "00001001101111010111110000101101",
602 => "00001111100111101110100010001110",
603 => "00000011011101101000100111001010",
604 => "11110011010011100110110100010110",
605 => "11110001110011101100110110001110",
606 => "00000000101100101010101001000010",
607 => "00001110110010000011011001100101",
608 => "00001011110010111110001011111000",
609 => "11111011001100000100111011101000",
610 => "11110000001000110000101010010001",
611 => "11110111011001110011100000011101",
612 => "11110011010011100110110100010110",
613 => "00000110000111110111100000110110",
614 => "00001111110111001111010101101111",
615 => "00000010000101101010001001101110",
616 => "11110001001101111100100110011011",
617 => "11110110010000101000001111010011",
618 => "00001001101111010111110000101101",
619 => "00001110110010000011011001100101",
620 => "11111101111010010101110110010010",
621 => "11110000001000110000101010010001",
622 => "11111001111000001000011111001010",
623 => "00001100101100011001001011101010",
624 => "00001100101100011001001011101010",
625 => "11111001111000001000011111001010",
626 => "11110000001000110000101010010001",
627 => "11111101111010010101110110010010",
628 => "00001110110010000011011001100101",
629 => "00001001101111010111110000101101",
630 => "11110100001101000001110100001000",
631 => "00001001101111010111110000101101",
632 => "00001101011111101000011110010000",
633 => "11111000100111001010110100010101",
634 => "11110001001101111100100110011011",
635 => "00000100110011111011000100011000",
636 => "00001111100111101110100010001110",
637 => "11111101111010010101110110010010",
638 => "11110000000000111110011000111111",
639 => "11111111010011010101010110111110",
640 => "00001111110111001111010101101111",
641 => "00000011011101101000100111001010",
642 => "11110000101111011001001100111110",
643 => "11111001111000001000011111001010",
644 => "00001110001100010011001001110010",
645 => "00001000100110001100011111100011",
646 => "11110011010011100110110100010110",
647 => "11110101001100001100100010001010");
begin

    main : process(address_cos_0)
    begin
        dout_cos_0 <= my_Rom(to_integer(unsigned(address_cos_0)));
    end process main;

end Behavioral;

