----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/18/2023 07:33:48 AM
-- Design Name: 
-- Module Name: cos_rom_1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cos_rom_1 is
    generic (
	       WIDTH : integer := 32;
	       WIDTH_2 : integer := 64;
	       WIDTH_3 : integer := 96; 
	       WADDR   : integer := 8
    );
    port(
        address_cos_1 : in  std_logic_vector(WADDR-1 downto 0);
        dout_cos_1    : out std_logic_vector(WIDTH-1 downto 0)
    );
end cos_rom_1;

architecture Behavioral of cos_rom_1 is
  type mem is array ( 0 to 215) of std_logic_vector(WIDTH-1 downto 0);
  constant my_Rom : mem := (
  
0 =>   "00001001101111010111110000101101",
1 =>   "11110001001101111100100110011011",
2 =>   "11111101111010010101110110010010",
3 =>   "00001111110111001111010101101111",
4 =>   "11111001111000001000011111001010",
5 =>   "11110011010011100110110100010110",
6 =>   "00000110000111110111100000110110",
7 =>   "11110001001101111100100110011011",
8 =>   "00001110110010000011011001100101",
9 =>   "11111001111000001000011111001010",
10 =>  "11111001111000001000011111001010",
11 =>  "00001110110010000011011001100101",
12 =>  "00000010000101101010001001101110",
13 =>  "11111001111000001000011111001010",
14 =>  "00001001101111010111110000101101",
15 =>  "11110011010011100110110100010110",
16 =>  "00001110110010000011011001100101",
17 =>  "11110000001000110000101010010001",
18 =>  "11111101111010010101110110010010",
19 =>  "00000110000111110111100000110110",
20 =>  "11110110010000101000001111010011",
21 =>  "00001100101100011001001011101010",
22 =>  "11110001001101111100100110011011",
23 =>  "00001111110111001111010101101111",
24 =>  "11111001111000001000011111001010",
25 =>  "00001110110010000011011001100101",
26 =>  "11110001001101111100100110011011",
27 =>  "00000110000111110111100000110110",
28 =>  "00000110000111110111100000110110",
29 =>  "11110001001101111100100110011011",
30 =>  "11110110010000101000001111010011",
31 =>  "00001110110010000011011001100101",
32 =>  "00000010000101101010001001101110",
33 =>  "11110000001000110000101010010001",
34 =>  "00000110000111110111100000110110",
35 =>  "00001100101100011001001011101010",
36 =>  "11110011010011100110110100010110",
37 =>  "00000110000111110111100000110110",
38 =>  "00001111110111001111010101101111",
39 =>  "00000010000101101010001001101110",
40 =>  "11110001001101111100100110011011",
41 =>  "11110110010000101000001111010011",
42 =>  "11110001001101111100100110011011",
43 =>  "11111001111000001000011111001010",
44 =>  "00000110000111110111100000110110",
45 =>  "00001110110010000011011001100101",
46 =>  "00001110110010000011011001100101",
47 =>  "00000110000111110111100000110110",
48 =>  "11110000001000110000101010010001",
49 =>  "11110001001101111100100110011011",
50 =>  "11110011010011100110110100010110",
51 =>  "11110110010000101000001111010011",
52 =>  "11111001111000001000011111001010",
53 =>  "11111101111010010101110110010010",
54 =>  "11110000001000110000101010010001",
55 =>  "11110001001101111100100110011011",
56 =>  "11110011010011100110110100010110",
57 =>  "11110110010000101000001111010011",
58 =>  "11111001111000001000011111001010",
59 =>  "11111101111010010101110110010010",
60 =>  "11110001001101111100100110011011",
61 =>  "11111001111000001000011111001010",
62 =>  "00000110000111110111100000110110",
63 =>  "00001110110010000011011001100101",
64 =>  "00001110110010000011011001100101",
65 =>  "00000110000111110111100000110110",
66 =>  "11110011010011100110110100010110",
67 =>  "00000110000111110111100000110110",
68 =>  "00001111110111001111010101101111",
69 =>  "00000010000101101010001001101110",
70 =>  "11110001001101111100100110011011",
71 =>  "11110110010000101000001111010011",
72 =>  "00001001101111010111110000101101",
73 =>  "11110001001101111100100110011011",
74 =>  "11111101111010010101110110010010",
75 =>  "00001111110111001111010101101111",
76 =>  "11111001111000001000011111001010",
77 =>  "11110011010011100110110100010110",
78 =>  "00000110000111110111100000110110",
79 =>  "11110001001101111100100110011011",
80 =>  "00001110110010000011011001100101",
81 =>  "11111001111000001000011111001010",
82 =>  "11111001111000001000011111001010",
83 =>  "00001110110010000011011001100101",
84 =>  "00000010000101101010001001101110",
85 =>  "11111001111000001000011111001010",
86 =>  "00001001101111010111110000101101",
87 =>  "11110011010011100110110100010110",
88 =>  "00001110110010000011011001100101",
89 =>  "11110000001000110000101010010001",
90 =>  "11111101111010010101110110010010",
91 =>  "00000110000111110111100000110110",
92 =>  "11110110010000101000001111010011",
93 =>  "00001100101100011001001011101010",
94 =>  "11110001001101111100100110011011",
95 =>  "00001111110111001111010101101111",
96 =>  "11111001111000001000011111001010",
97 =>  "00001110110010000011011001100101",
98 =>  "11110001001101111100100110011011",
99 =>  "00000110000111110111100000110110",
100 => "00000110000111110111100000110110",
101 => "11110001001101111100100110011011",
102 => "11110110010000101000001111010011",
103 => "00001110110010000011011001100101",
104 => "00000010000101101010001001101110",
105 => "11110000001000110000101010010001",
106 => "00000110000111110111100000110110",
107 => "00001100101100011001001011101010",
108 => "11110011010011100110110100010110",
109 => "00000110000111110111100000110110",
110 => "00001111110111001111010101101111",
111 => "00000010000101101010001001101110",
112 => "11110001001101111100100110011011",
113 => "11110110010000101000001111010011",
114 => "11110001001101111100100110011011",
115 => "11111001111000001000011111001010",
116 => "00000110000111110111100000110110",
117 => "00001110110010000011011001100101",
118 => "00001110110010000011011001100101",
119 => "00000110000111110111100000110110",
120 => "11110000001000110000101010010001",
121 => "11110001001101111100100110011011",
122 => "11110011010011100110110100010110",
123 => "11110110010000101000001111010011",
124 => "11111001111000001000011111001010",
125 => "11111101111010010101110110010010",
126 => "11110000001000110000101010010001",
127 => "11110001001101111100100110011011",
128 => "11110011010011100110110100010110",
129 => "11110110010000101000001111010011",
130 => "11111001111000001000011111001010",
131 => "11111101111010010101110110010010",
132 => "11110001001101111100100110011011",
133 => "11111001111000001000011111001010",
134 => "00000110000111110111100000110110",
135 => "00001110110010000011011001100101",
136 => "00001110110010000011011001100101",
137 => "00000110000111110111100000110110",
138 => "11110011010011100110110100010110",
139 => "00000110000111110111100000110110",
140 => "00001111110111001111010101101111",
141 => "00000010000101101010001001101110",
142 => "11110001001101111100100110011011",
143 => "11110110010000101000001111010011",
144 => "00001001101111010111110000101101",
145 => "11110001001101111100100110011011",
146 => "11111101111010010101110110010010",
147 => "00001111110111001111010101101111",
148 => "11111001111000001000011111001010",
149 => "11110011010011100110110100010110",
150 => "00000110000111110111100000110110",
151 => "11110001001101111100100110011011",
152 => "00001110110010000011011001100101",
153 => "11111001111000001000011111001010",
154 => "11111001111000001000011111001010",
155 => "00001110110010000011011001100101",
156 => "00000010000101101010001001101110",
157 => "11111001111000001000011111001010",
158 => "00001001101111010111110000101101",
159 => "11110011010011100110110100010110",
160 => "00001110110010000011011001100101",
161 => "11110000001000110000101010010001",
162 => "11111101111010010101110110010010",
163 => "00000110000111110111100000110110",
164 => "11110110010000101000001111010011",
165 => "00001100101100011001001011101010",
166 => "11110001001101111100100110011011",
167 => "00001111110111001111010101101111",
168 => "11111001111000001000011111001010",
169 => "00001110110010000011011001100101",
170 => "11110001001101111100100110011011",
171 => "00000110000111110111100000110110",
172 => "00000110000111110111100000110110",
173 => "11110001001101111100100110011011",
174 => "11110110010000101000001111010011",
175 => "00001110110010000011011001100101",
176 => "00000010000101101010001001101110",
177 => "11110000001000110000101010010001",
178 => "00000110000111110111100000110110",
179 => "00001100101100011001001011101010",
180 => "11110011010011100110110100010110",
181 => "00000110000111110111100000110110",
182 => "00001111110111001111010101101111",
183 => "00000010000101101010001001101110",
184 => "11110001001101111100100110011011",
185 => "11110110010000101000001111010011",
186 => "11110001001101111100100110011011",
187 => "11111001111000001000011111001010",
188 => "00000110000111110111100000110110",
189 => "00001110110010000011011001100101",
190 => "00001110110010000011011001100101",
191 => "00000110000111110111100000110110",
192 => "11110000001000110000101010010001",
193 => "11110001001101111100100110011011",
194 => "11110011010011100110110100010110",
195 => "11110110010000101000001111010011",
196 => "11111001111000001000011111001010",
197 => "11111101111010010101110110010010",
198 => "11110000001000110000101010010001",
199 => "11110001001101111100100110011011",
200 => "11110011010011100110110100010110",
201 => "11110110010000101000001111010011",
202 => "11111001111000001000011111001010",
203 => "11111101111010010101110110010010",
204 => "11110001001101111100100110011011",
205 => "11111001111000001000011111001010",
206 => "00000110000111110111100000110110",
207 => "00001110110010000011011001100101",
208 => "00001110110010000011011001100101",
209 => "00000110000111110111100000110110",
210 => "11110011010011100110110100010110",
211 => "00000110000111110111100000110110",
212 => "00001111110111001111010101101111",
213 => "00000010000101101010001001101110",
214 => "11110001001101111100100110011011",
215 => "11110110010000101000001111010011");
begin

    main : process(address_cos_1)
    begin
        dout_cos_1 <= my_Rom(to_integer(unsigned(address_cos_1)));
    end process main;

end Behavioral;


